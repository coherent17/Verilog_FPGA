module piano(rst,pb,clk,seg0,seg1,seg2,seg3,seg4,seg5,one,two,three,four,five,six,led,segh,segt,sw);
	input pb,clk,rst,sw;
	output one,two,three,four,five,six,seg0,seg1,seg2,seg3,seg4,seg5;
	output [9:0]led;
	output [5:0]segh,segt;
	reg seg0,seg1,seg2,seg3,seg4,seg5,clk1,clk2,one,two,three,four,five,six;
	reg [4:0]state,nstate;
	reg [23:0]count,count2,i;
	reg [6:0]ledstate,nledstate;
	reg [9:0]led;
	reg [5:0]segh,segt;
	//frenquency division and change the clk1 is a function of t 
	always@(posedge clk or negedge rst)begin
		if(~rst)begin
			count=0;
			clk1=0;
			i=0;
		end
		else if(count==5000000-i&&count>=1000000)begin
			count=0;
			clk1=~clk1;
			i=i+25000;//every period the count will minus 100000 so that the frequency of the clk1 will increase
		end
		else if(5000000-i<1000000) i=4000000; //the speed wouldn't become unlimit at last
		else count<=count+1;
	end
	//debounce the pushbotton
	debounce o1(.pb(pb),.clk(clk),.npb(npb));
	/*always@(posedge clk or negedge rst)begin
		if(~rst)begin
			count2=0;
			clk2=0;
		end
		else if(count2==(5000000-i)*2)begin
			count2=0;
			clk2=~clk2;
		end
		else count2<=count2+1;
	end*/
	//memory logic for the segment state
	always@(posedge clk1 or negedge rst)begin
		if(~rst) state=0;
		else state=nstate;
	end
	//nextstate logic for the segment state
	always@(state)begin
		if(state==5'b11111) nstate=5'b0;
		else nstate=state+1;
	end
	//output logic for the segment state
	always@(state)begin
		case(state)
			5'b00000:begin
				seg5=0;
				seg4=1;
				seg3=1;
				seg2=1;
				seg1=1;
				seg0=1;
				segh=6'b011111;
				segt=6'b011111;
			end
			5'b00001:begin
				seg5=1;
				seg4=0;
				seg3=1;
				seg2=1;
				seg1=1;
				seg0=1;
				segh=6'b101111;
				segt=6'b101111;
			end
			5'b00010:begin
				seg5=1;
				seg4=1;
				seg3=0;
				seg2=1;
				seg1=1;
				seg0=1;
				segh=6'b110111;
				segt=6'b110111;
			end
			5'b00011:begin
				seg5=1;
				seg4=1;
				seg3=1;
				seg2=0;
				seg1=1;
				seg0=1;
				segh=6'b111011;
				segt=6'b111011;
			end
			5'b00100:begin
				seg5=1;
				seg4=1;
				seg3=1;
				seg2=1;
				seg1=0;
				seg0=1;
				segh=6'b111101;
				segt=6'b111101;
			end
			5'b00101:begin
				seg5=1;
				seg4=1;
				seg3=1;
				seg2=1;
				seg1=1;
				seg0=0;
				segh=6'b111110;
				segt=6'b111110;
			end
			5'b00110:begin
				seg5=0;
				seg4=1;
				seg3=1;
				seg2=1;
				seg1=1;
				seg0=1;
				segh=6'b011111;
				segt=6'b011111;
			end
			5'b00111:begin
				seg5=1;
				seg4=0;
				seg3=1;
				seg2=1;
				seg1=1;
				seg0=1;
				segh=6'b101111;
				segt=6'b101111;
			end
			5'b01000:begin
				seg5=0;
				seg4=1;
				seg3=0;
				seg2=1;
				seg1=1;
				seg0=1;
				segh=6'b010111;
				segt=6'b010111;
			end
			5'b01001:begin
				seg5=0;
				seg4=0;
				seg3=1;
				seg2=0;
				seg1=1;
				seg0=1;
				segh=6'b001011;
				segt=6'b001011;
			end
			5'b01010:begin
				seg5=1;
				seg4=0;
				seg3=0;
				seg2=1;
				seg1=0;
				seg0=1;
				segh=6'b100101;
				segt=6'b100101;
			end
			5'b01011:begin
				seg5=0;
				seg4=1;
				seg3=0;
				seg2=0;
				seg1=1;
				seg0=0;
				segh=6'b010010;
				segt=6'b010010;
			end
			5'b01100:begin
				seg5=0;
				seg4=0;
				seg3=1;
				seg2=0;
				seg1=0;
				seg0=1;
				segh=6'b001001;
				segt=6'b001001;
			end
			5'b01101:begin
				seg5=1;
				seg4=0;
				seg3=0;
				seg2=1;
				seg1=0;
				seg0=0;
				segh=6'b100100;
				segt=6'b100100;
			end
			5'b01110:begin
				seg5=1;
				seg4=1;
				seg3=0;
				seg2=0;
				seg1=1;
				seg0=0;
				segh=6'b110010;
				segt=6'b110010;
			end
			5'b01111:begin
				seg5=0;
				seg4=1;
				seg3=1;
				seg2=0;
				seg1=0;
				seg0=1;
				segh=6'b011001;
				segt=6'b011001;
			end
			5'b10000:begin
				seg5=0;
				seg4=0;
				seg3=1;
				seg2=1;
				seg1=0;
				seg0=0;
				segh=6'b001100;
				segt=6'b001100;
			end
			5'b10001:begin
				seg5=0;
				seg4=0;
				seg3=0;
				seg2=1;
				seg1=1;
				seg0=0;
				segh=6'b000110;
				segt=6'b000110;
			end
			5'b10010:begin
				seg5=1;
				seg4=0;
				seg3=0;
				seg2=0;
				seg1=1;
				seg0=1;
				segh=6'b100011;
				segt=6'b100011;
			end
			5'b10011:begin
				seg5=0;
				seg4=1;
				seg3=0;
				seg2=0;
				seg1=0;
				seg0=1;
				segh=6'b010001;
				segt=6'b010001;
			end
			5'b10100:begin
				seg5=1;
				seg4=0;
				seg3=1;
				seg2=0;
				seg1=0;
				seg0=0;
				segh=6'b101000;
				segt=6'b101000;
			end
			5'b10101:begin
				seg5=0;
				seg4=1;
				seg3=0;
				seg2=1;
				seg1=0;
				seg0=0;
				segh=6'b010100;
				segt=6'b010100;
			end
			5'b10110:begin
				seg5=0;
				seg4=0;
				seg3=1;
				seg2=0;
				seg1=1;
				seg0=0;
				segh=6'b001010;
				segt=6'b001010;
			end
			5'b10111:begin
				seg5=1;
				seg4=0;
				seg3=0;
				seg2=1;
				seg1=0;
				seg0=1;
				segh=6'b100101;
				segt=6'b100101;
			end
			5'b11000:begin
				seg5=0;
				seg4=1;
				seg3=0;
				seg2=0;
				seg1=1;
				seg0=0;
				segh=6'b010010;
				segt=6'b010010;
			end
			5'b11001:begin
				seg5=0;
				seg4=0;
				seg3=1;
				seg2=0;
				seg1=0;
				seg0=1;
				segh=6'b001001;
				segt=6'b001001;
			end
			5'b11010:begin
				seg5=1;
				seg4=0;
				seg3=0;
				seg2=1;
				seg1=0;
				seg0=0;
				segh=6'b100100;
				segt=6'b100100;
			end
			5'b11011:begin
				seg5=1;
				seg4=1;
				seg3=0;
				seg2=0;
				seg1=1;
				seg0=0;
				segh=6'b110010;
				segt=6'b110010;
			end
			5'b11100:begin
				seg5=1;
				seg4=1;
				seg3=1;
				seg2=0;
				seg1=0;
				seg0=1;
				segh=6'b111001;
				segt=6'b111001;
			end
			5'b11101:begin
				seg5=1;
				seg4=1;
				seg3=1;
				seg2=1;
				seg1=0;
				seg0=0;
				segh=6'b111100;
				segt=6'b111100;
			end
			5'b11110:begin
				seg5=1;
				seg4=1;
				seg3=1;
				seg2=1;
				seg1=1;
				seg0=0;
				segh=6'b111110;
				segt=6'b111110;
			end
			default:begin
				seg5=1;
				seg4=1;
				seg3=1;
				seg2=1;
				seg1=1;
				seg0=1;
				segh=6'b111111;
				segt=6'b111111;
			end
		endcase
	end
	//memory logic for ledstate
	always@(negedge rst or negedge clk1)begin
		if(~rst) ledstate=0;
		else ledstate=nledstate;
	end
	//nextstate logic for ledstate
	always@(negedge clk or negedge rst)begin
		if(~rst) nledstate=0;
		else if(ledstate==7'b1000101) nledstate=7'b0;
		else if(seg0==0&&npb==0) nledstate=ledstate+1;
		else if(ledstate>0&&seg0==1&&npb==0) nledstate=ledstate-1; //no light but push 
		//else if(clk1==1&&ledstate>0&&seg0==0&&npb==1) nledstate=ledstate-1; //have light but don't push
		
	end
	
	//output logic for ledstate
	always@(ledstate)begin
		case(ledstate)
			7'b0000000:begin
				led=10'b0000000000;
				one=1;
				two=1;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0000001:begin
				led=10'b0000000001;
				one=1;
				two=1;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0000010:begin
				led=10'b0000000011;
				one=1;
				two=1;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0000011:begin
				led=10'b0000000111;
				one=1;
				two=1;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0000100:begin
				led=10'b0000001111;
				one=1;
				two=1;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0000101:begin
				led=10'b0000011111;
				one=1;
				two=1;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0000110:begin
				led=10'b0000111111;
				one=1;
				two=1;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0000111:begin
				led=10'b0001111111;
				one=1;
				two=1;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0001000:begin
				led=10'b0011111111;
				one=1;
				two=1;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0001001:begin
				led=10'b0111111111;
				one=1;
				two=1;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0001010:begin
				led=10'b0000000000;
				one=0;
				two=1;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0001011:begin
				led=10'b0000000001;
				one=0;
				two=1;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0001100:begin
				led=10'b0000000011;
				one=0;
				two=1;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0001101:begin
				led=10'b0000000111;
				one=0;
				two=1;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0001110:begin
				led=10'b0000001111;
				one=0;
				two=1;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0001111:begin
				led=10'b0000011111;
				one=0;
				two=1;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0010000:begin
				led=10'b0000111111;
				one=0;
				two=1;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0010001:begin
				led=10'b0001111111;
				one=0;
				two=1;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0010010:begin
				led=10'b0011111111;
				one=0;
				two=1;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0010011:begin
				led=10'b0111111111;
				one=0;
				two=1;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0010100:begin
				led=10'b0000000000;
				one=1;
				two=0;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0010101:begin
				led=10'b0000000001;
				one=1;
				two=0;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0010110:begin
				led=10'b0000000011;
				one=1;
				two=0;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0010111:begin
				led=10'b0000000111;
				one=1;
				two=0;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0011000:begin
				led=10'b0000001111;
				one=1;
				two=0;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0011001:begin
				led=10'b0000011111;
				one=1;
				two=0;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0011010:begin
				led=10'b0000111111;
				one=1;
				two=0;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0011011:begin
				led=10'b0001111111;
				one=1;
				two=0;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0011100:begin
				led=10'b0011111111;
				one=1;
				two=0;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0011101:begin
				led=10'b0111111111;
				one=1;
				two=0;
				three=1;
				four=1;
				five=1;
				six=1;
			end
			7'b0011110:begin
				led=10'b0000000000;
				one=1;
				two=1;
				three=0;
				four=1;
				five=1;
				six=1;
			end
			7'b0011111:begin
				led=10'b0000000001;
				one=1;
				two=1;
				three=0;
				four=1;
				five=1;
				six=1;
			end
			7'b0100000:begin
				led=10'b0000000011;
				one=1;
				two=1;
				three=0;
				four=1;
				five=1;
				six=1;
			end
			7'b0100001:begin
				led=10'b0000000111;
				one=1;
				two=1;
				three=0;
				four=1;
				five=1;
				six=1;
			end
			7'b0100010:begin
				led=10'b0000001111;
				one=1;
				two=1;
				three=0;
				four=1;
				five=1;
				six=1;
			end
			7'b0100011:begin
				led=10'b0000011111;
				one=1;
				two=1;
				three=0;
				four=1;
				five=1;
				six=1;
			end
			7'b0100100:begin
				led=10'b0000111111;
				one=1;
				two=1;
				three=0;
				four=1;
				five=1;
				six=1;
			end
			7'b0100101:begin
				led=10'b0001111111;
				one=1;
				two=1;
				three=0;
				four=1;
				five=1;
				six=1;
			end
			7'b0100110:begin
				led=10'b0011111111;
				one=1;
				two=1;
				three=0;
				four=1;
				five=1;
				six=1;
			end
			7'b0100111:begin
				led=10'b0111111111;
				one=1;
				two=1;
				three=0;
				four=1;
				five=1;
				six=1;
			end
			7'b0101000:begin
				led=10'b0000000000;
				one=1;
				two=1;
				three=1;
				four=0;
				five=1;
				six=1;
			end
			7'b0101001:begin
				led=10'b0000000001;
				one=1;
				two=1;
				three=1;
				four=0;
				five=1;
				six=1;
			end
			7'b0101010:begin
				led=10'b0000000011;
				one=1;
				two=1;
				three=1;
				four=0;
				five=1;
				six=1;
			end
			7'b0101011:begin
				led=10'b0000000111;
				one=1;
				two=1;
				three=1;
				four=0;
				five=1;
				six=1;
			end
			7'b0101100:begin
				led=10'b0000001111;
				one=1;
				two=1;
				three=1;
				four=0;
				five=1;
				six=1;
			end
			7'b0101101:begin
				led=10'b0000011111;
				one=1;
				two=1;
				three=1;
				four=0;
				five=1;
				six=1;
			end
			7'b0101110:begin
				led=10'b0000111111;
				one=1;
				two=1;
				three=1;
				four=0;
				five=1;
				six=1;
			end
			7'b0101111:begin
				led=10'b0001111111;
				one=1;
				two=1;
				three=1;
				four=0;
				five=1;
				six=1;
			end
			7'b0110000:begin
				led=10'b0011111111;
				one=1;
				two=1;
				three=1;
				four=0;
				five=1;
				six=1;
			end
			7'b0110001:begin
				led=10'b0111111111;
				one=1;
				two=1;
				three=1;
				four=0;
				five=1;
				six=1;
			end
			7'b0110010:begin
				led=10'b0000000000;
				one=1;
				two=1;
				three=1;
				four=1;
				five=0;
				six=1;
			end
			7'b0110011:begin
				led=10'b0000000001;
				one=1;
				two=1;
				three=1;
				four=1;
				five=0;
				six=1;
			end
			7'b0110100:begin
				led=10'b0000000011;
				one=1;
				two=1;
				three=1;
				four=1;
				five=0;
				six=1;
			end
			7'b0110101:begin
				led=10'b0000000111;
				one=1;
				two=1;
				three=1;
				four=1;
				five=0;
				six=1;
			end
			7'b0110110:begin
				led=10'b0000001111;
				one=1;
				two=1;
				three=1;
				four=1;
				five=0;
				six=1;
			end
			7'b0110111:begin
				led=10'b0000011111;
				one=1;
				two=1;
				three=1;
				four=1;
				five=0;
				six=1;
			end
			7'b0111000:begin
				led=10'b0000111111;
				one=1;
				two=1;
				three=1;
				four=1;
				five=0;
				six=1;
			end
			7'b0111001:begin
				led=10'b0001111111;
				one=1;
				two=1;
				three=1;
				four=1;
				five=0;
				six=1;
			end
			7'b0111010:begin
				led=10'b0011111111;
				one=1;
				two=1;
				three=1;
				four=1;
				five=0;
				six=1;
			end
			7'b0111011:begin
				led=10'b0111111111;
				one=1;
				two=1;
				three=1;
				four=1;
				five=0;
				six=1;
			end
			7'b0111100:begin
				led=10'b0000000000;
				one=1;
				two=1;
				three=1;
				four=1;
				five=1;
				six=0;
			end
			7'b0111101:begin
				led=10'b0000000001;
				one=1;
				two=1;
				three=1;
				four=1;
				five=1;
				six=0;
			end
			7'b0111110:begin
				led=10'b0000000011;
				one=1;
				two=1;
				three=1;
				four=1;
				five=1;
				six=0;
			end
			7'b0111111:begin
				led=10'b0000000111;
				one=1;
				two=1;
				three=1;
				four=1;
				five=1;
				six=0;
			end
			7'b1000000:begin
				led=10'b0000001111;
				one=1;
				two=1;
				three=1;
				four=1;
				five=1;
				six=0;
			end
			7'b1000001:begin
				led=10'b0000011111;
				one=1;
				two=1;
				three=1;
				four=1;
				five=1;
				six=0;
			end
			7'b1000010:begin
				led=10'b0000111111;
				one=1;
				two=1;
				three=1;
				four=1;
				five=1;
				six=0;
			end
			7'b1000011:begin
				led=10'b0001111111;
				one=1;
				two=1;
				three=1;
				four=1;
				five=1;
				six=0;
			end
			7'b1000100:begin
				led=10'b0011111111;
				one=1;
				two=1;
				three=1;
				four=1;
				five=1;
				six=0;
			end
			default:begin
				led=10'b0111111111;
				one=1;
				two=1;
				three=1;
				four=1;
				five=1;
				six=0;
			end
		endcase
	end
endmodule

module debounce(pb,clk,npb);
	input pb,clk;
	output npb;
	reg [2:0]shift_reg;
	always@(posedge clk)begin
	shift_reg[2:1]<=shift_reg[1:0];
	shift_reg[0]<=pb;
	end
	assign npb=(shift_reg==3'b110)?0:1;
endmodule
