module shiny(led,clk,rst,sega,segb,segc,segd,sege,segf);
	input clk,rst;
	output [9:0]led;
	output [7:0]sega,segb,segc,segd,sege,segf;
	reg clk1;
	reg[9:0]led;
	reg[22:0]count;
	reg[4:0]state,nstate;
	reg[7:0]sega,segb,segc,segd,sege,segf;
	//reduce the frequency
	//original clk run 2500000times get the inverse clk1;
	//so the clk1 T=2500000*2=5000000 get 2Hz clk1
	always@(posedge clk or negedge rst)begin
		if(rst==1'b0)begin
			count=0;
			clk1=0;
		end
		else if(count==2500000)begin
			count=0;
			clk1=~clk1;
		end
		else count=count+1;
	end
	//memorylogic
	always@(posedge clk1 or negedge rst)begin
		if(rst==1'b0)state=0;
		else state=nstate;
	end
	//next state logic
	always@(state)begin
		if(state==5'd29)nstate=4'b0000;
		else nstate=state+1;
	end
	//output logic
	always@(state)begin
		case(state)
			5'b00000:led=10'b1010101010;
			5'b00001:led=10'b0101010101;
			5'b00010:led=10'b1010101010;
			5'b00011:led=10'b0101010101;
			5'b00100:led=10'b1010101010;
			5'b00101:led=10'b0101010101;
			5'b00110:led=10'b0000000000;
			5'b00111:led=10'b1000000001;
			5'b01000:led=10'b1100000011;
			5'b01001:led=10'b1110000111;
			5'b01010:led=10'b1111001111;
			5'b01011:led=10'b1111111111;
			5'b01100:led=10'b0111111110;
			5'b01101:led=10'b0011111100;
			5'b01110:led=10'b0001111000;
			5'b01111:led=10'b0000110000;
			5'b10000:led=10'b0000000000;
			5'b10001:led=10'b1000000000;
			5'b10010:led=10'b1100000000;
			5'b10011:led=10'b1110000000;
			5'b10100:led=10'b1111000000;
			5'b10101:led=10'b1111100000;
			5'b10110:led=10'b1111110000;
			5'b10111:led=10'b1111111000;
			5'b11000:led=10'b1111111100;
			5'b11001:led=10'b1111111110;
			5'b11010:led=10'b1010101010;
			5'b11011:led=10'b0101010101;
			5'b11100:led=10'b1010101010;
			5'b11101:led=10'b0101010101;
		endcase
		case(state)
			5'b00000:sega=8'b11111110;
			5'b00001:sega=8'b11111101;
			5'b00010:sega=8'b11111011;
			5'b00011:sega=8'b11110111;
			5'b00100:sega=8'b11101111;
			5'b00101:sega=8'b11011111;
			5'b00110:sega=8'b11111110;
			5'b00111:sega=8'b11111101;
			5'b01000:sega=8'b11111011;
			5'b01001:sega=8'b11110111;
			5'b01010:sega=8'b11101111;
			5'b01011:sega=8'b11011111;
			5'b01100:sega=8'b11111110;
			5'b01101:sega=8'b11111101;
			5'b01110:sega=8'b11111011;
			5'b01111:sega=8'b11110111;
			5'b10000:sega=8'b11101111;
			5'b10001:sega=8'b11011111;
			5'b10010:sega=8'b11111110;
			5'b10011:sega=8'b11111101;
			5'b10100:sega=8'b11111011;
			5'b10101:sega=8'b11110111;
			5'b10110:sega=8'b11101111;
			5'b10111:sega=8'b11011111;
			5'b11000:sega=8'b11111110;
			5'b11001:sega=8'b11111101;
			5'b11010:sega=8'b11111011;
			5'b11011:sega=8'b11110111;
			5'b11100:sega=8'b11101111;
			5'b11101:sega=8'b11011111;
		endcase
		case(state)
			5'b00000:segb=8'b11111101;
			5'b00001:segb=8'b11111011;
			5'b00010:segb=8'b11110111;
			5'b00011:segb=8'b11101111;
			5'b00100:segb=8'b11011111;
			5'b00101:segb=8'b11111110;
			5'b00110:segb=8'b11111101;
			5'b00111:segb=8'b11111011;
			5'b01000:segb=8'b11110111;
			5'b01001:segb=8'b11101111;
			5'b01010:segb=8'b11011111;
			5'b01011:segb=8'b11111110;
			5'b01100:segb=8'b11111101;
			5'b01101:segb=8'b11111011;
			5'b01110:segb=8'b11110111;
			5'b01111:segb=8'b11101111;
			5'b10000:segb=8'b11011111;
			5'b10001:segb=8'b11111110;
			5'b10010:segb=8'b11111101;
			5'b10011:segb=8'b11111011;
			5'b10100:segb=8'b11110111;
			5'b10101:segb=8'b11101111;
			5'b10110:segb=8'b11011111;
			5'b10111:segb=8'b11111110;
			5'b11000:segb=8'b11111101;
			5'b11001:segb=8'b11111011;
			5'b11010:segb=8'b11110111;
			5'b11011:segb=8'b11101111;
			5'b11100:segb=8'b11011111;
			5'b11101:segb=8'b11111110;
		endcase
		case(state)
			5'b00000:segc=8'b11111011;
			5'b00001:segc=8'b11110111;
			5'b00010:segc=8'b11101111;
			5'b00011:segc=8'b11011111;
			5'b00100:segc=8'b11111110;
			5'b00101:segc=8'b11111101;
			5'b00110:segc=8'b11111011;
			5'b00111:segc=8'b11110111;
			5'b01000:segc=8'b11101111;
			5'b01001:segc=8'b11011111;
			5'b01010:segc=8'b11111110;
			5'b01011:segc=8'b11111101;
			5'b01100:segc=8'b11111011;
			5'b01101:segc=8'b11110111;
			5'b01110:segc=8'b11101111;
			5'b01111:segc=8'b11011111;
			5'b10000:segc=8'b11111110;
			5'b10001:segc=8'b11111101;
			5'b10010:segc=8'b11111011;
			5'b10011:segc=8'b11110111;
			5'b10100:segc=8'b11101111;
			5'b10101:segc=8'b11011111;
			5'b10110:segc=8'b11111110;
			5'b10111:segc=8'b11111101;
			5'b11000:segc=8'b11111011;
			5'b11001:segc=8'b11110111;
			5'b11010:segc=8'b11101111;
			5'b11011:segc=8'b11011111;
			5'b11100:segc=8'b11111110;
			5'b11101:segc=8'b11111101;
		endcase
		case(state)
			5'b00000:segd=8'b11110111;
			5'b00001:segd=8'b11101111;
			5'b00010:segd=8'b11011111;
			5'b00011:segd=8'b11111110;
			5'b00100:segd=8'b11111101;
			5'b00101:segd=8'b11111011;
			5'b00110:segd=8'b11110111;
			5'b00111:segd=8'b11101111;
			5'b01000:segd=8'b11011111;
			5'b01001:segd=8'b11111110;
			5'b01010:segd=8'b11111101;
			5'b01011:segd=8'b11111011;
			5'b01100:segd=8'b11110111;
			5'b01101:segd=8'b11101111;
			5'b01110:segd=8'b11011111;
			5'b01111:segd=8'b11111110;
			5'b10000:segd=8'b11111101;
			5'b10001:segd=8'b11111011;
			5'b10010:segd=8'b11110111;
			5'b10011:segd=8'b11101111;
			5'b10100:segd=8'b11011111;
			5'b10101:segd=8'b11111110;
			5'b10110:segd=8'b11111101;
			5'b10111:segd=8'b11111011;
			5'b11000:segd=8'b11110111;
			5'b11001:segd=8'b11101111;
			5'b11010:segd=8'b11011111;
			5'b11011:segd=8'b11111110;
			5'b11100:segd=8'b11111101;
			5'b11101:segd=8'b11111011;
		endcase
		case(state)
			5'b00000:sege=8'b11101111;
			5'b00001:sege=8'b11011111;
			5'b00010:sege=8'b11111110;
			5'b00011:sege=8'b11111101;
			5'b00100:sege=8'b11111011;
			5'b00101:sege=8'b11110111;
			5'b00110:sege=8'b11101111;
			5'b00111:sege=8'b11011111;
			5'b01000:sege=8'b11111110;
			5'b01001:sege=8'b11111101;
			5'b01010:sege=8'b11111011;
			5'b01011:sege=8'b11110111;
			5'b01100:sege=8'b11101111;
			5'b01101:sege=8'b11011111;
			5'b01110:sege=8'b11111110;
			5'b01111:sege=8'b11111101;
			5'b10000:sege=8'b11111011;
			5'b10001:sege=8'b11110111;
			5'b10010:sege=8'b11101111;
			5'b10011:sege=8'b11011111;
			5'b10100:sege=8'b11111110;
			5'b10101:sege=8'b11111101;
			5'b10110:sege=8'b11111011;
			5'b10111:sege=8'b11110111;
			5'b11000:sege=8'b11101111;
			5'b11001:sege=8'b11011111;
			5'b11010:sege=8'b11111110;
			5'b11011:sege=8'b11111101;
			5'b11100:sege=8'b11111011;
			5'b11101:sege=8'b11110111;
		endcase
		case(state)
			5'b00000:segf=8'b11011111;
			5'b00001:segf=8'b11111110;
			5'b00010:segf=8'b11111101;
			5'b00011:segf=8'b11111011;
			5'b00100:segf=8'b11110111;
			5'b00101:segf=8'b11101111;
			5'b00110:segf=8'b11011111;
			5'b00111:segf=8'b11111110;
			5'b01000:segf=8'b11111101;
			5'b01001:segf=8'b11111011;
			5'b01010:segf=8'b11110111;
			5'b01011:segf=8'b11101111;
			5'b01100:segf=8'b11011111;
			5'b01101:segf=8'b11111110;
			5'b01110:segf=8'b11111101;
			5'b01111:segf=8'b11111011;
			5'b10000:segf=8'b11110111;
			5'b10001:segf=8'b11101111;
			5'b10010:segf=8'b11011111;
			5'b10011:segf=8'b11111110;
			5'b10100:segf=8'b11111101;
			5'b10101:segf=8'b11111011;
			5'b10110:segf=8'b11110111;
			5'b10111:segf=8'b11101111;
			5'b11000:segf=8'b11011111;
			5'b11001:segf=8'b11111110;
			5'b11010:segf=8'b11111101;
			5'b11011:segf=8'b11111011;
			5'b11100:segf=8'b11110111;
			5'b11101:segf=8'b11101111;
		endcase
	end

endmodule
	