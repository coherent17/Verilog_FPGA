module ictexampleseven(a,o);
	input a;
	output o;
	assign o=~a;
endmodule
